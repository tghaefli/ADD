XlxV62EB    6431     ca0Q+�d���&�Y|\k��8���x��K�.v03��{���>R�F�#�Q5*� ����q��[�8�-pd7��.��{f����|j诂i���'c3q��H��4=a�Ŝ<l�L��J�n���X(��Y����[��|�Vh�0���Ь�ʭ�=H�vC��ڀz?�ԏ{qK

X
"=%�"�#����9����Q��P�aFjQ��`�GϮ�+䘮�dm5�
f�&mQA��<xxl�6=�V����Ҩל������[�Zv����4�%b��_�[UU`ܣ��!�`ܢ�$s�y�ek�W�L��l`K.";c�?��6�Q�>�yL�R��&�+�����i�u��z:�(z.�p��1<�Αz�î����j���L�J�q�ܿ{�䅲���sD���Y��g�V�p��^�W�F�a����$ԗ�,��M���Ȕ�t\�U�ǩ&���[sM��4�.�6���R!�/��f���������НG��D1t��i>n�G�^7��r�{����� n�y����H%�7K��<����ĳ��I�ʬ�q�^�y����(�:�n\�C7&��-|�q�]��?�p!�P��>�N>O��D��o�1aF�ɫ���f���j�&��̘���@S�|�r�ftS�&aj�U���5<���v��{U��S͡󧆽��;���w�SA�+�zU:�T[5C��m|aq'w�c tw�EE�����is=��.����nD�=C���5�9#��v�5:}G�v�d7ک��}�y��˅��_d�P��	W"*��E#���d��1p��8*WHW}�B�0D}�R�u�(-pr��asc��V�nR=�]�4>�@�����D<Z`�e�A�$�?J��Ӯ:H �xS�-2Q0t�Cʶ)2�[[��aqMd��kUh�� ��gIN%���֊�%�j-�ر\|P��i���9�R� G��j�6%%g0�J����@�I�Sui�Αpއ&�YE��O�sǄ�i�zF��y�VՋ+�-�$�"�&���H@�,+깽��gN��*"�Y�~ܾQ2"'�3 ׯ�ui��J�3v&��\R5������~����N��������p��N|��1%j���^(�Ŀ9�Z��L���[� �����֖�l��	Ӟ�n�4�+����	v�:�"�sfϹ��c^b���\��U3�c�G���lӱK���[�M������!(EGFԍL�\�����B���Ec+����O��s���K�^��bQBP������<Z����e�t%HY�\���.0z��}^I {εYSO�z��'���O�3�*{����%'���,RI��B�z��Na�_ʶJ���ǫ�<?��j#[���4�:yUf���E���=���u��[�˨�E��|�>G����e��4������Z8��ӂG�^t͹Qo���*z���[�������(T�=��Vkc[���ԅL�?�>�2��*���1=��SK/;3��ץT�=Q�:�8Z��/�C����*X�c�I��R�����q����������Mo5���*�s<�I���!"P>��e�����v�Xç���q�@��g�������u�jƯ�S�I1=k?��P��.�Q4K�#Ȍ5����<_أ����Gd��!Ͼ��Y��.x�ǚ����kYܜf�|�Hg,�ܕu0�yq&N����oZ���1���V�dP��.�4��E4FP$E���x �6zd{�q��s��J�T��W��u�ʣ;����~RW|�>��l)+@>U�)
�ty]U|�;ݖ���l���d}�s��Z��TU�$��'�0�[j�+x�͆�����Ck0�j�����)	+��$�s�#�ϮiO�Ӵ �і��yJ�C��TI���̔!t+�QT3H�����˺�����Z�2�0�q1��o6�&3��-W��b��D����������G�Z2k!��Ͷ����i����`�k�2*4 ��+e�Oh�KA�XG;^��⫈���ƫ'��D�?���͇�P6���f�������/��5�*6t�L���;`c�a܎��q�ˣ�����=4~5$�T�KӉ]��S8�� ��(=Tm��1�6��8m-H�%<��i���Fw'�S�\TB����w ��J���a��)��r�����z:}��5-��{�.�����0�(�R���VD�q�:���HI��%�$�P�Zf�����omu���BL&�&њ���F��Hnc�N9-�ʨ���q���e�i�j��GGe�A����Xx�X�3�l�4�?�|;��Qf^)�p�Ӷu��wޯQ��7H[�Щk�O�i`�(F�a��~o@J��F�_"�ٺgk8�YMp�$��^)�p�bZ���B�@�9"ySF
5��'8����2T�ׁU��r<v�`�Q�_U�B���_�"�Ι�S�hN�4��G��k2WCF�-\R8-Q��u�жu+Ym�ލ����Y��Ѿ��n��!�}f�&��+�,�(����y�Z#�D�i���᝖;�ft��I �){6��g��4Mj퇼�[�-T��	#vq׍��g�o0Lqg�c��T�1�w[��C�S��z�ag�a�+k$)"����@�����)�8�������+�E�&��ww��މ2�6�R�jҬq�<ٌ_���]{ZFNf��W��UA�˄j^��-hܰ�q��8��.��>�]SO(M��ޮ+Ju��ϒκ%ES�Q�>Z^�NG�)g2a�-��+ {�~w��P�볓=Υ�Z���s�����l���K��:��?l�;�����W���W:��~Ԛ��RW�}'�3yi���4�l>a�$��+E-����q�!���'1	�3�*����h ;�H�Մ͕-5��/Ň��fB�5�*C��ߍ �U��/~x�7ʕ���T��3*���Z�#�8��4��Ѭ�����Sg��)�&����ү@aq�;+FM�b>�g��/�K�A�Xg�8����G��7c�==�?d��?f_n��>�(���������O�jj���A�UTc,��ѿ�7��"��x��B��v��'�P\�����&��D�cP�T|`.��x�!�V٫(8�-C�3�̳G`F:����}�Y�����c��:�,��(2��3�8��L�p��sg�h,�Z���<��	1Z.