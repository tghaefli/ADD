XlxV62EB     754     240�Z)H��2�k��*	���a��ƞ�� -��ü�����ܯ� 2�V�*��P�=S���cu��L4�	蒭ЄIś�N�v�����F����&]*ETx���U��U�Ы��:�E�� pk���\<��6V����<z[�T�|�=	�K��#+��JL�5��5���s+ߥn���ڱ�^� a�N���ۈ���`����@��J�j����q>ۅ��!ya��9����O�v��W��Ҝ��@ۨ����h�eB�T~�궷5���B�n��c<p�� G��Y`��-:�=��#��G{v�M0Kx���:��ñ�d^��^�����e�t��W��e��I��>Q�!�����yd��m*��ٱ�}Ga ��wi��mB������~'j��$��a�}^un���sQ�� �"��ھ'��ǱV��&YP�y�!�0'K�A���E���@Hw�A�R�v��<֦��;u@q�[��j��
a��z����	�&���u1˯`FK�pu��<�t(��\��$���]a������������I�D��<��͖�h�F�
�����ʹ�PaU/