XlxV62EB    fa00    22d0�x���u	�]*��D7�������Dln���Ԋ��{�h$*Ϥl<�LE�/���7Ŝr	�R�Ub}2½}���sqj�7@��<z�{����"�n�>�������卻b�:-�3��?a�M. �ڣ�@��i�"�WHP��c �ΝH��#�����l���R���h�}�L2�Y�W��ku�N���#�������EP6Q� �(���؄�����X�߮�cǆ��Z�����9?�8<�Ǟ���F�$�t9X��g��N��e�T��U�d
 �.��4*��sG�/�rP��#m�`y�&�#��D�z�u��0���s��`h���t@�]�Y`�%�Tw��$�9��{�)JM�ON�"�����#��7xc����d� 
rO���-H��q�[q�[�j�>�&�s>�S��G��CÍXd4�. �,��ʴ�:�T��?e	����~��~ʻ��P'3g���e\���/k�J��� lo����;C|�0v���UZI7#�bl�p�#X_���?�ɾ����>�'T�G�D[���Ŗ�7x��v:��o��<��
 ́���S�1����BU�3��N�L6y0��^i��/d��]���	r1w�;�	�΃F�h���O�)\z;Mf�>�7��l+�}�4���73�87��XHp,���c%��Y0$�I��z6�}g����,�2'���^�4��a�N�YE����2�C�lo{�j�MH�?0�|��L�滎�D?If�;S!�zX��F� I�P`-��� ����������^���\���5(�&�DR�-��l1h�@��Q�yB������%B�yv�
��'cc�s��mO�m`�v����gi忧��������q��z�0��:N��x7SC`p2����և�TjXq:�J�C-������]������\� E�{���iI���]�AU
�r�tA��ϐN�r7cFpQ�c^�#��Kb�W����b�/�+v?�� ),H/��I���D���b|���E�Y@s��W���q���g��r������e��<pD�߱��L����-2W���M~��-Jq �Z�~�Ċ�Am��㖔�i�;�������rϪG����7�������nRմ���*G��ê�T(���7��JM��������_;O�7Lm(�w�Q��r~����n�n�eU�+�A�BT���'�p�X0|;�B=68u���]�@M/�9
��K������/uYC��6*������ ���(�8��9:��ۜK�@��*��DNF�dyce��k_������N4J��[���F��)������yQ�k�.j߫5�L~�h�����~"��ECFs�jYbVѷ�Jmی'� ���6*�<xQG���-�iAЬ����o�������=��0�1��;g���^�,�MTp:8����(��ϥ��iC������N)OL�H�d%�zg��SG���[�O:�l]@�8`��W���d��PD�F������i������K�X��l�*�����
�(xT72�WH4�����B�=�<�6�D��k8�����W/0��9+/���5G y�S�]��������M焝��才4�a�U[A�~�N�bW]A�_���Pƴ#�̵��NG7x����ӯ�7��2⡎�����b���a-��U�gf7����AD�?�?a��"d�@M�G�*w�F:K���!8�&�P��w��Ğ�-�2nzNF��{�$b�5���ޮ���}� �1�!�z<�ʒK��������@��z���O;LL�#~ZXui��y9�q�fa/.J�3����Ł�w��\�^�)N����u�Z!?�^y�+�z_و{�Nv���6�(-������JqY�6}
�"�^��x�+	�/�琭X�3F(Ӟ؞��F
r ���R;Һ뢡KpQ~о,��V��p�e4��w�3������.<Z>r�jN�Xw?�:�?���T->��I�,�t*�0c!'!�_?��e���v�%�x��и诬v�wzN���5��,o�UK����.m0���}p�@b����o�-�(u�������6��O<!�BAS��4�8�T�"�H��5@_�u��0�<U��(�^ah�Mw��&�6��٣�6�ڸ�wd������1��!n���L�0Oz����HU��e_#�����'H��5���8�x�q᛬C�x��C��v�����_MJ_������-��O�5L�W�fK�s1[����+�&���d����_:���{������WzAf�����jg��	G������28�=՜��0ǟ�����d������"S$���{��*�Dt28������P\��@:�M*�IqDyPZM�H�sV�aUt^ڊ�Fa4rIuxC��(����+�5Z.���_FAĳ2�F�ʓ�vzY�s��H�2�%W�zB�;��+k�̷�E�9N ������T@���Ď.h\+r�mlÑ��1T먣����-�ȱʩp*<�'V�|����hNs]�7��M6�zt#����O#,��X֢��^��:����;6��D���>X3���� aT�l�>�%�IzO���dFqq��P3���������2T�a��Y�@$��e[7�EZQ���DT���7���̮2~H�o�Uc��,�ߕ�.`O�7jU�5r�xR��~%q���3���"q��+b���.���?B�R���Z��<_�!�Z���v���H������(���ݫnk�sc}(x��՝F��H�?<iƟ�&����y%ФUt�S�RR�>�q*+�E �O���*2���ֲpc5ƫ��[�mbA}@lS'@��`�ec�����s�Y���M.�>:%��@݃�s�GɄ-�R7�y�삇�8l��<���d���i��p�Jb����/o�F�%g&�nZ�
�*xA��tiO�(8̈��"v4��i�2�g�4XCFCQ����C�Q7?����9�:~�V���Gɲ��K��b���Y6��� ��bJ,��'��)p��ы�Ex����'���I��_�j{�(|�*�u���������L��Y��S1�]��9��k�m���9�',�XO�:Lv�5��J��]@����p���N}hjf�	��c�~T�B��°Ci�HE�ˤ�[S5�/�Ƽ�c=Ԙ�#2Q�3`㮧Ri�1ѧ0���"+�	���\η�~3�Ձ\CFᘆV ��C�_[xH)�6��*?����SԸ:�$U���R�\&4���.wӆ0�M4O�h<�M#�����b�Exǆ }SW���v2�RW��[i�7&�7������o���'"�n1)�U�'UB��hyy�@ņ�$�բ�Gǉ� C�&�����y}���<�f� ����v4�'
�*K��k@��X�x�p�L�;���h81M�j�
�|�@,����n��R�~��a�~��L㷐�G��VX�M�712=����Nf%�u�<��|~-� 杠vܙ�}0��B+��8��2���;�/%�;z�wk�DU�y^6��4�_������(ƫ"�7=��F�-"�*��S���C_N�PY���W�v�R�(|�����`6�L�:�LZ�&!)}�Lp����Z텰�o��Cr5���Ȗ'�730����#�����T-=�f�����UQ����V���"n
��F�[�N���\2���{���y�S	�DBڐ�r.���`"�b)��9`�<'�n��|;�4Zx�hNr�1$dHu�_�U�q>�1�޼��U�����9ʮ�'6��n��3�f�-5�}L��$���0τ��R�t��A�b��p�Y�Q+ ��=�9X�)���{�˘@ʁzɺ�B�J&�|t� ��d"��tr���h�B�ˠ�(V�fr�Be��0\��C_����6k1!����N�.5�:C�Rt��O>Jd�ŔH�M"�~�O��%�P��"�*����هa׎����������{���5�p�x#��l����v�SP%z������5�ZzE��.�6ˠ3�� 5�$�yk�!�
^�3;�)��[+N��$��D������B�]�nκ�&����6E�y��e>b_����.� ⵡ����(f,��^AXy��`~��e�l�k� s��$�`����J!���/���m#��r��W�].ϝeC��������P���緀 ��H�-튨�]��҅@3��Ժ���F4蘿6
�5/Q$OӄD�h8��Y��\*R���L@z�s�R35 .$��Ы�L, �o�������E�����wr���H��QY��@���F��,���.���> �I�4��^�.d����4SBp�i��O�֜���@�I��G)���ED�/z�%b��o���Y6Y`{�a��3*�ғx�s^�H`&;@�]�3��=����0 �y� �YoS��d&l:��H���ۘV2��_�+�D"���z��p�8���tܧ�\9���<б���u���dв3mY�P[\ J�'���,�v�Y.6��O0 WJ�zi��:	L����n� �`&����R��n��堭�_��Ōo����<`=}Sa�8�����#V����(���|]LEn���a�F�:H9��d_n~Cu��-$���ۈ��ٵ,M;��)����Ep"C��&�n���_����O�tv����Q�RSM^���C�_}�T$�B��s��@����G�Y0��H4��g�9W�\��L'yf���k��ٽXQ�Ћ!��z⡣}�|��A�b�X98�e�i��,�2W:��h�.�e�������U~��Uw�0�J����嚿G4��b�Z�	����{�ƽ[�aV�	�|R�@��ɬ͌{��V�7Z��}�{(8p�>��p�%��~y�π�h ��ol��K��#�w ���v�/�T炫ܐ�|k��/����� ��N�}F[d@isҒ�ΰߢPN�?C:�F���R{�J�+�Z�&���C��-��eP^|�P#��vhu�!�y�3�;a0e1�W�Ӯ�*%�K+4�	�MK0��{�1D�a�T>��Z(��'hC� :V�S��&���}�R����C��
��+�
_6�z/���T8�S��L��2���?���2V��w���0��B��[՘���Q���/3��N��.�HT�Z��I�yd���^ϸ�������>�4����Dʷ��U[�ėg"}g>�X�`�lx��$Я���n�	"�����m����6TV:B��������dP`�@ ߁�dY��^j_�8����sw$hT�{L���~�p���������(�Z�+����[1��j�]�!�HTI��cK�9���'��ear',�`�cY�a
x�:�L5�V��S��(�ɂ!�q;Zge�q~�<W(&����VC[�����Z�O 2���)=7^*�Qs��Z�?����1��g��	��1��@�=�N����<��#|	����v����ٌ[Zh�\r�װ����` �
�O�]� ~9�W ��+�ô1�R�w�k�="�Y�f���J��g�{�)}f�P�Ä�Փ)��֟����b��6��;H�[>�U�0�`Ft�H�!�2��#4�%�7T[QK��.�X4N#u�`�꽱�҅-���~�~�͛%����5]��M�PÆ��K��[A�L���ؘp��t���ԉ�%������,���X�ye%w���{*_�Q��23��Ԧ���D�F�k�+L�0�h�`{R�)��,zɣY�ր�#"R)���˚���w:�?���,�E%���])Y�%��ߋH*�Y,�>�=�l�O���+��R,g��	�睕��ܦ.6ͅ�Μ�~��>��d�f[� ����-`�+Cnxޜ��˧B�\�,�/ο'5�ZX�謚��v|��Y`�m�W����L�*�ٱC�ݝ��R
B��M�b^�p��߰�AE<����^��DWge�3�i���ۑ�&W�;#�����^��le�6��ώ�'�6���?��5���Ǵ6tQ���4�zy�-]SGD��f�>�G�׋���uf�Q�1n@c��cn�)2�En��¾��r���0Q&r�m	�U������3��S��^9f�2�f�J�L�&Y$Jq{���.pы�5�mo|L�P�6��n�݆p#��+|9/�0�2J%�3|ᒱ8����ω�ئ�lUofU`Mґs�e�GC�X9^�ZdHS�#	'�:]����o����L���ۋg�㴸o�<U��R:��q����h��픩ƍ�e��,׎�=^����?���(���N%���W`���b��Hb:JMզ�]�8�G��l�~��5�׎�E�ơ��- �l���R_�#
u�hm��M��}�w�lv��u���l������ն��M� '�/��}t�9����4�RC5)=jQى��9�[��6C�͑G\8!؅Oz �Q������[~��˔JX�Fp����=�s1D��8b�M�>ߵ��"���|7��`Fa��K&XXq�CRi/����W+�
�P�����錶9�Br5��z�/���o��]dQl�i�}?���O��a����a���jL!��`�<�������(�b��ͻ1���]M������ɗ=i.f����w?qp��3n�B�3��c%�Ƅ��2��6�����){��b\���l��c�x"�O�sNF�J��Xs���Z�������l�w����(XG�%��$*&��B���!'N�n��{�z~�"��=I$�-��Hf����lƷuC$5u��wH|�զ�C�%����]By\����g[��8C�@�}��Oj�䊁�`Q��Zq=!�@��M;&1�D�D�VԌ�Ss��p�oW�w&w�J���⍩�hL�}�'��q(��N���K�����ҍV�)�Ҙ[t�v7*�J��U��j���w��CwK��u�H�$��HF������:oC��qy�������b����Y4�k�i�/l�N���%ۥ�B�(#��K�ϱD܎�._�aa��>i�oa�%P�^R��YfE�Ϛ�d�A�HnW�vN�ό�p��,�5�����~K%�y}�#�m(r!m�y;iS-6V޿��3v�*w��s�h1/�
f���N��5��2w��2�d��6��m��)z����U�A���VC��"�2D����4�甡9��H��O��"#�s_yy��N��
a=� ��ED���M�5��Ῠn�l�\efJ8�_=;�j��!��|�Xy��Ex�A�T+�X/0�^'������%�3�Y�5b���ށlޕ*4��18���C���K��v��Z�	T�*Z���/tUHF�)��?v��~�ܵ�?�����3�p�q-cu\aV&j7/�w+��g��J�>fiB_d��\h~y�g�	Bȅ�p�6T��@�S� !V�A%V��?�p:��ϻ´)������u�@E���w�2Ji
��Sf s��ԗo��<X>�<O圩f��i,����.n^P�/�qG��qy�+��e:���\f�|~"-�� �)�Rcar�p�ڪ��y�����HiA�pr�o�K����֧S��ڢ]�����! �<^�Z��C;���(�g�o	�0�:3��ྠd�,�a/B��`����<.�e�jf���s[��1r��..ÓM+���@o(7P��\�s9N���=9h�U�S�8���k�"�(��'����zTi�A�d���+���a��,�lX��3@��W㗹��A�����t���������4P��4����p�/c{�QOK��Ҩ=M~3���c�̐��Q~haK�B�ߋg�Fh6�7���N�d�:�� �����PFF�ls��"�A��,A��%\����z�/�*�P'�Q ��5����CQ��C#o&N�2�V5z���'CH�-Ȳ��L�*�Br������J�5���22u{��>�/m�D�Hl]��=�!^���܄�G�dIAd���t��b�������:Eu�D\�U��&���k�A"f~^�?f�
�z;EM8���w����FA�2C�n"���ĮmZn���n���H3>mU�=�t��>��#��������,�v4�R����R��4���9#.R=�-Ϡ75�[/��9]Wd�֓.�fE	���� ;F�.���-.O$��#�
 �	�i���_�
H�#��IT�Ɓ����j�0���Rz�*�`"��DUp��7���7�³qd��%d��U�P���ޑN�ݗ�/��6��8���m����	c���I���v��[Tr�%xG�
%SEk��@�� �)e:so��a����`�p�U�	|�,;Ym���ͣ�B��!��I�b*�(a��m�޷����c�c�b�9ڠ�q���c��=�Q���'�q�*;~�v9r_�Ϥd��+xb;���X-I+b�*���Q@�!�\Q�n2[����rl�5�#jL�]��3���j���R�V�
��.�B���7C���o?uD�_K_J�b\�6�*Աxy1��BY�C��lEo�v�l��ZW�&�Y6�>�pJ��TE�M�i(j�!_�E.N�R��_8�S��j��Е:)--�IG[b�{�%�<���Hcr2�*;�)�'���lA��Wh l��iicS쿋Ig?,�j�1��Ч�g�m4�+���Ⱦc��\(�Z���9�}�nJn�.XlxV62EB    4c04     900��S�v�k->C@����o��c`�8�IHl����5�l��ߙP��b>A�
h9�Y[D=HF������j�8f�R�L�Kb]e�v�K�`�9�HS;gL[ن�
����2�;��ׅ���[�r��V��LMH����3E٨p>�F��7\�V�p����Y��S�zAJ�a8~�l��nR���'�9%�,��l!�׋b��}~?L`����?X��[JK�T�M��(�U�*Ag�XH6CjƟ:�C��%/���l0U����F����~��_�)	��	Irb�]ɖ&��o����_�Y\��:����EBR�`�6&��Y��?2Pٰ�9�u���yu$-i�m`�/9z֩�fx�
r棶��TQٟ枀�����jd�H�//�,����lRcLzZ--��n��DofTYI���)s���D5�����1��=�_��_5��N�8�k����eR��X�!.���W�,#�蘟�1���k#pa���޼������K��ɻ��=)�����i�'3C/�G��/a*�m*li�x�$��^1Z�%���	ﺍ.P�U���&h{noY�Ի�f�*������6T^�-�wN��ՏJ6\�Tkj��	tԭ͠�|�#l?��N�w�.��@��PJ�PNi��n^E18O�̯:ܿ3# �8w����[9�8�fi����w�k  �R��Mr�ұ�Z�x ��
"%i�։�	ڿ��a,?���FY�Pl)��:J��\ "[���t�/m�ImJs	�[u4�.�GXկW̗RsV��������Ծ�ޮn�0�|Y����6�0�T��ۀ�I�T4$s��v[0��?Xp���n������i���l�J��g�׀�9�˻�(l|.�
e�i����Q:�׏�tF��0T�"���ú,�D�,���K ��zC�n���m�EUA�M�F�
��|C�>Z�S��QF5�M���e�D�f��w�=<\�Hq��m�cb�\���\2�\�3��fͪ#$L
{f����R�������ct!�7z:c�`��!�� 9�X��t��5@i���¿M�9M�Vi���_m^�H������j�{#`,���;��\&�MS�x��>��'a�H�����d�v1�I�i U���gZ�����3m�N�kw���E)/�Me�>� 
�	a�߾KEz�A�9H(>3ŵ�)�(���
K>�Q��a�˿�0���,HY���A{��uQ�R�"q��~�Z4��Ѡ�&� ���813l}%��?�Q=���Pj_���v�?Y�v�=_�����V�;��L.��š���	4�C��d�
$	N������@�=�ILA�T�W�2߃����XU��P�UR�*�S̥EQ�9e'�Q�		�Dj����J@�.P/�T�����ȯ����qIt(Wl8��;��t@�r�lb��N��q��5}���?�0<�q��-6܍l���=n�F�Vh)��3��!�% ����H��b�d]���b<�W8r�JY�Y������;��>8v̓˛��T[Ep�t\<-,˕*��zѻ�
�8��aGMJ>�_5li���섦DS�`k%�텎��O���;��Dx�����m˴��D�H�IJ��(�e�P
���+��\{��Wm9��~k���],�������}\Lܕū�O�����{K�LF�[4��l��K?�����_a!��k����7�C�a�U�Zm�}{��^ⴟ���\W���Bsno9$�A
�S����N��wK���+���z˃{'p^�CcQf�W,%R��?9��c�CQ�G�X4L�n��)���Ϯ)���_/���e��"�6��է�h/C��)�{�+�<��jR%�-�t�C�@��o^�u4�hM�SB��o�N�w�6U�󸣺qf{i��?(��u �$v��ٴM3���t7;��lP�PW�{%�����sD���[}-��s��U{Tf �����X��a��\q�_��E��t�Љ!��,f�n΍":B�֤eJ���ݐQ�6���xF�L��H��x1���&U[/���y4jl"��S�B��@QB��������P�$' I:��呢�fo���Sm;�O�>�&f������Z�?��\�<��8ʸ�h���A��0a�̞�Ŕ��E�v��.��T�fR�IɁ~�Sf^�X������39�C���+SI��s�r	T�V��zV4D3��	�Kz"��<��=��\NT���w�P(>wtw�	k�,X=����