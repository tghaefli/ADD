XlxV62EB    2245     e00W��[K���,��2u�.*��bV<�>铓�Ԏ�%w���]5@y��qZ�,�{3蹮SU�f���ߊ'8���T������!ǔ�q�M���&b3������+�{����y��2n�Zg'b�s�D�M*��粞�Щ��
�͈�;ș�rUh�3�j0O[&�_�x��%ӧ��"&����m���NO$8~4HP�����i�SNM�d1�|�3�L!�*�Wx`L8��]A��<��g���o��ۿ},�O����`�x�Ng-o��_�ȍR���TIA412�����^��-��U�F�J��R5p!��^�$g&�n�z��T)ԉ��d�'U2Pܵ9��j�I��D���jQ(�K���X6�����v]�:	��+m���Og�< &6٦�������������b�3�\x����1V,������C?\R�7K����$�6��������
��$r d�A�szm����ޟ�����y���N��Ar���i"?c�WN7W��G�Z��,�dP���Lª������B�������Y�+gN���ʈ�U!v(��#���&m��Gh.���:�+2�=���F}6�?�8�r����4%�5(Iq��(m�Dn�E�dX��v�%(�
*�}�k�����6j|",��I�q'�<���"�"܂>͉y�T	n�B�R�����/����3nՒ6d�g~ 9\��ת���_1���hh)jg��\���)p��CL� ��*�$x��>�z�ܘ�Z�k7����x2����z��e�(��<G�~�]G�A��\�� *�D��p�-�S&��y��I��I�2�g>�>�������z����/�J*�� ��=��x�m|«���4n�v�i�������ʬf��jRn��tgKع{'�)bQ�˺a��� ;�K���u�?�3r�- �V������$��3�����Y]?$=���si���Ŕ�w��A��7�s������b��5Dް�aO��]����^Pn��V2�Ah������ro�c�����\�0��6�oQ�NŻ���gR	.R��Z�zǄ��:�ȣ�;O�h��R�Y%�1��:�,W�WF��<J�cb�O����������y2�����!�=Ӌ-܇�d72���)Є�>g�Mo'_M�{��##���7���K ����r�H�4qG���`��G[2�[�ؕy��G�y�/���ڤ�"�kT`�KB͸%�!6�=�!6����j��2�caC�j�P������3Z +��H����"�֔�l|�u�@ ���ȂT�D8�{��$��d�2�NsփM��l�5_�%�[�j�53e]�������k(dm8����^}��
��oT�/_�M}���2�r�r�t�n����gwջ���a"^�u��7�P�ȫ�[�b�XB1���.W�$�����>kD��az�a1���O�D���vi�J$�h� J}�����u�0�uW��:}�)����7��/{���1,#Y"p�$���R_osvq1%����B߯}���JB�_Ȩ3Mmﱣ�d�^�f��;�������Y���٣�Ɯb���ߊ����Ԡ��ŵ���Y��8��zQROs�N��P�ڷ?����q��J��t�y��ϴ����܆hB�Qh�i������O]����?.< ���2+RjpH����өҽ�aN@�2�~��f�--��s@�Q�L�Lr��#;�F��ೇS*�U�G�ot�V�O����Õ���oҩ �"��P�F*פ���4�@Jx��s���`���aW���ײ8VOJ�Q��q�7�~q�Tؒ��]�|���
�f�ToFFNR*Ǯ@����чoVSb��V����o嘭߇��d�[�Y�v~q����u���γ��*ylH�{a�d� 3A��ܾ�Sb�=��č4�V��\n�9@�@[�]N��ꪩP�����1���	���?�ou�AkZtQ`��Q�<�=h�5-���b2ٚF�o?y����r(��բpLXc�~����"+��2��(�繑0����s�]n��å��txFӱ>�Dh����o�K�ɺHe�|H�s�oDa3
o5�׫����zQ%���͌�xro���b�Ǝ��[�F��ȏ�������u�H���Y�K�ӑ��G�.����B	������>͵��D����;��3���aD~{��J�>����y�uM�36J��]J��ԇ�/$ �Za4.�!����<]y{.'�:��:����'v�,����1_���������13|-����K�Q:��1u\=��D�::���mpԃ""2��F֫�.�o!㺢J�O�+�V��)�B4�Zc�����I=�lr:v%`�nRp	$H+��%Gjj��$h2�x���7�V�IJ��'���z�/<.F�Ӕ����&�6����Hx9�f�jl���=&�Г��ъ��oM;�P�=aĈ�7}�W.B�˝\�ڋ��v�e��ሯ�e���F�����ȃ�C��!��7�H��'�jLӫs��8��]a���^�=8���������J*�\�Ft�Us��Z.3Lf�x+�x��W����y��kݭ��[���T]��?XNWS�m�.9l��inPY�_����g �	OX.Di&:�B,���=޾��d��⟫ՍY�XaQ��:���O'��0B�{��@�q��^	`��Q��#�>��қL�f��#\a<��-(�)�
[���TXE�qs+:�9�:l��*�C �����N�����Ҁ*nS� �6ּ�oF�2�XB=��K����n�*�)���5�7T���`�$��s�/�s�~d�\9����T�n&�[���v����r�����z$c���Z�|������[�p*�4�Ș�&W�q�7laX��#/n�Эq�$&��?�6�p�x�y2��Co����C`����s܋�M�*�_>�m��6vx��mh�ť�攅F��@[�V fC �^f(�����>}֊�c�e�p���)ƅ�k�����D��)|�K�i�c�z]/.6���>�����b6BI ����A�;�+7��K����=(���;���ٴ�璢��@��&~ymj���~v��R,"ػ�sK�	2T�^���G�g�Bp�kËq^@*1��V���|�Rn?��������n���G^P�ԑ�w�/��\s H���¿t�V��	�lb̳Zǆ�5�l:�HI�d�Zp����Zp�3���BS9
 ��~;>c`/�<�c��3����s��G/33�C��t/�$��|S�/�=k�L[�߆��f7]8���x�12�:�c�)��Bir�сLVA��� ?!58l�a�l(Y�L�+�B�E��!�hߔ�Z��l�W��84?��Q�W�/NA^1L����6B�Yu���t)l�?���UI���L���z�Բ 軩�*�λ||�U<�a�q�.tE͹?.�=���wy<\����o�܃��o��t�S��r_�