XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$��^�M5o�j�bӗ��満{[�	��7�2��'�i.�ܰ�T�W��N�fj���v�`Z���ï]K����`~ȃ)n'�7���	-�%e*�n[L���#x���I.Z���%�����Z���H�� uv&P"�͋mxL�@@e�&EO5QަG�\�^�h`{�{"��e�\���ř,�=EYp&XǑV[뼓�!�_�gBS�P/*�a�i��41o�w��:�9�a�o�s�J�]�%s��mI*��qS��M�]ﭞ4�r0?n�T�sT�}���Ίa~j�5�z�ς������#	�$p�'J���8�z�G�St<�Q@v#~B
H��P5d��g��=U�MqoG��i�e|Jц���^|�Kl�˅Q��V
��k�s>��<Q�}�2�@���Q #{�g ���\�x��M��2�
��>�#A�n���f'�K�-�6j�SR���?2��� ��$�(s�g�,�#��R�'�J~�`{�p>�Gus�E{=)t�1���T{��*���n��ق��(�E�a��Q���zouU�f��y��lU��5UB��BA\�mF��f��}�N[<FUxy���� S�v!����͓ɸ"�N�}^��}g���2H1}�v5���ܕ�*�i��T���Jyx �U�3����J7�r���7��/dC"�X���a�R�sl�Xe�m�l���2<#y��'31Bl����1���!�=�W%���\{��l�	$[�C?XlxVHYEB     400     170�^m�c�5��&�T��~���T��������?I�S۸�-\S���XTd*.�yz�e)b��$������1ﳫ����j�<>,�f��o������ c�\pu��~�|7Oy�i�y�����҃�UvxBZ���x�����G0�0�m�/�5�9o�x�h��Rf	}qԜq���ssɌS��l���k�U.�W�Kx��n��.�/� \�~0(Ԉq��l�4�$� �y��F�	l>7� �� SH(>�^3��\��2H��e����P,W��
w9�j ��|Yς�S�n�|_k7+�#���Z��vh��3g��,M`R�ZΤ�Y����1�<M�TH�/N���H+l)YW2��6"XlxVHYEB     400     1b0'�Fs���W$��Ry�!�[�_`����|��5���s9'�=Z��:՚p�u��K
�7�v����p�+Kg3�f���~��-y��Q�/8~3��%�}�V���~�����\\�͂ۤ��KG�P�'C��=ReH�W���+:{�Eg��
	U�����K���&2���p����a!}-��r>3�3��o����&�z�e�r�oT��~����ߦóz�N���ژ6C�0nvȎh�y�����IK p��_��Y�e�� !����a�,A����ɲK��:Jr����� <}�|�������5�'���W��ڙ�N�L��L�[ŎL�Q����6��"�q�0Ur�]�wԙ9��瓩D��{��U����}��&�/g� ��z��a�ܪ(z=Y�p�w��g�'�J�mj�,XlxVHYEB     400     170�.R����M�>����C��d��������y�TugM8VDR
_ɑU�{;E��r᭐f�e٤�@�P;h�C�*2]��Im�	E�2�����ct=Gz˝���E���R& �4q��X��_I�ؼ`/W���\����Ge�	밴,���\��RH��}�5���V幗��Q�`���2�Jj��Rl���r@d�l�p��Vbo��/��y�����l)�۞��W^���
wbK�yjH�`�8�$QY_�bjF
�{�d��s��G���*��
��qI���6����ն�C��O����.��[��]^nEeX�Tz�YDu��h�?G���?�:aB�Ě_ɿ��:5[��9N�XlxVHYEB     400     170�_�GPP)<@�Y��髽�
���]q�ρv�y+��Ta��l����1�/8���2A+�_��P�r��Z����e�F�~��eB� �]|��m�zH�.=���/�i���STj%�5�8�$4�y(�� �7���S�ψ�ۓ�@�=���/��xd2���^tFL�	�m��ߙU?��0	B�p�X�mr�S�<���,YxZ� �+xyϦ8��3,�ʶ~�čΔ$���,�$�)+q���h动鯽dAh�?�<6HC2�-�ԡ4��r�V�A�"	�m}8E	�����$i:1����U� 
�.@�5���:�F�Q�IG5�,P|>���͸&�A��^vXTreC����\ǭ�X�.�㏨�ڝ�R�`"YXlxVHYEB     400     180��Y�a�.�
y�~S�z��+JWQlk���]�y��R��&p�Fc����1/�M�	p^Je����/�Q9g:l��8r��K���`�j����:Ę�������h����(����ev���dχ���oQ������)�9�;�C Q�3`�yvb�tB7`�C+pj�I�D=W�4i�SM�1���2$ٜF7Y�'4Ԣ�n�NA��s|$�	Pl ۊn��_39�� ��Ї&��I�s1	��$N�j·Z;��k�چCzO����}��훹� �6|ܟ��4�ܜ�E�≑	�sE�K���ʭ-z�h����S@#��R�%3ؐUf����>��1�� ��~ٝ��@�n>���0�^��G����E��-�GXlxVHYEB     400     190�.M5����b?��mD ���-���wH)��N�n38~)����d	6�O����d�c��(v�D���/���hh�3����5Mcc������W�(���̆�	��a��=�$Qv{�����Ծ�)�3�!{�'�M�m�|�y��f����&s� ȷ%P��Dl߅��=?��Pl�\�A6L6�c�7͏v�R�t�b٫�*Ps�\Q��u~�$";n)�}R"�
�wL�iF�Ez��Th����A�S���fX�l=��|��1Ķ���"���׃���1{��1c�^u}�ҹ��9���G��%��Yښ��u6��|ओ�a��x@g���X����`, �΋��G���U��;�h.\�:�vhQ�t�Z�pj��@�^��XlxVHYEB     400     120��j�=�$(S���u���2|-�D�1Ū�����2Nc'��;��}�\ؖ���ᡧalۯ�Le?�B_�$�V]y�}�;�fb�����@���5�	ɨZ���d	�m���-��x���VcD�=�u�ꌟOxD�@kT���I]���Ɣ�z��'�W�F��Îxi% �qH>/Z	Fl��m��Z�%:]q�M��F��k:(ȥ҈�[�F-�?������
���{�%��9;��V�b2 �n�&T=�`5t2�����rᐯ�mE�R&���$٭u���0]�>XlxVHYEB     400     120�M����)ͩ�G.����"���\��{eH���U��"��Ћ�����ρ��B9��+C����Js�M"4OTY�u�X�,Ǽ~�L,��򅥌��y��e���A���U1����
G*k}b�TK��.~���I���/��7���G���5�%��z㬿#�E�Qn�~�3�9��>���TN£쮎lx�v��(�I+�][�2�4H�������b���Ddv����]��������`ٗ�;!�\��w̠d��1�����Nh�[���$E���XlxVHYEB     400     100W���.w���}��	S����#3��'��}_��Mչ�L�]N�R��T��֬e���0���X��$�@�d�!'��}|!�>�"��R�{���)Gfϒ������ܾeP`�-Q�`�� ?�����O�v�}#Cɯ�"�.��,���4���D�T�޾:c[͓-a��V▇C>��$����<��ˋ%n1���g�.��`��� �O���ҕ`�� K��
�٘x4�C�z�T�z56���$XlxVHYEB     400     150�B���+�
�r�,c�ΔB�:f[�砟�~Ի���s[�v�xV6�>zݢUW���� ��a��5|#�:��ᰙ�s	�q��jf1��]f���TY��ya�0W��&[�E+@f:��'$��vZ'���̦�3
� ��9�uck":�N�G��D�R{_F�:>W��������R��T8B��v���(�? �6%��o-�4�����M[��v�#H�l��ҝ� �Д�o�a���h`�������x-0�Z��Hĝ���c6`�#{J�<�����|�԰�l�|͒�}}'+QX����`��ʖS��]�ű�{k��B	���s��[����ÁXlxVHYEB     400     120hI�I�9���P�P
��<��o��>�J���.��\~.]Y��n�������2�Cf���}͎�ڄދ�tqY7u6t����eL��%g��Ǩ���s���eH���"~�����pd�bjMX��?�6�'����d;��y����a��ϚjG�8��yd;���z������EcW��{$�y�a�\�|��Eҽ����ͼ�هlU� dfT��if<�yҭ�}CՓ�h �:����:�2�P��(�v]�%���ΥZ�Q��1����}'�_><�)��ޜh��4�XlxVHYEB     400     170�������+�Ґљ3��ծ T����-J�>��-�Lô�ۧR=�X,�6��9ղ�QEԷz���tU���>��=e����\&a�F�]��B�:�/lp ��$	-�p���F�T�я���:ir�ǝ<���qZ$�C�غ7�H����/�'h�+�WN��u=<���s�V�LK��7$�{����C�̢/9��^O��lrrR��&��A0K�MY���=.�Y����mŵ���<X߀˩����;��_�.df���fr���V��!!C�Gª�w�M�� f���5j�?b����I)$���˩��RoNiq��MQ��a��)�Q[P�Vy: J�+gǒ�a���
L�2�XlxVHYEB     400     160Do��rN|�*��߯�V����Z_ϊ�D��K�qca �?d�\!jf#�IF4R�����-Tg��G��74_��Z��,��A�g�Z+�o�̰7�rx@=fŤ��aktW�^����'� �_+�^�DEL���X��{�ɷR�/,� �3B�4����Ԓ[�T�ѽ#7��Q`�Z9�_�1$�%�GD���~)ڔ-?�k�J+���������0V!),�x����B�$�K�'��B�:����m�t~3ƀW�r��ǅJE�($D�BX��%⸘�\����@�%mn�y�KT�DnR^C1m�Y	ʟ��u������`�&�N[�|��N�XlxVHYEB     400      e0g�
�+X��wz�^|�;�R�mmN����.�w��0@�aAfj�_�-�/�Bʊ���j�GI�s�P�,ZY' �дŜ���	��:zZ��k|(z�A�_:��kS�I��`7sY���^�N�H�B�Wu�-��a��;���Z���',�2�f*��L��I�{�מ*q�������o����&�<q�p�-XFnڐ��:?ޱ���^XlxVHYEB     400      c0K��%@�sбz\l\����G�O1e�~D��俅t�E,��8�
�Nw��F5c�����9K_o�B��G�3ÚzP���[�@�T�h��"�|[�eX�(q%���h�p����Y�8d�� ��!=Pu(��y۟eE[A�e�\᧬��)B����g�[����K�@5gt _�Q6������,�AQC&EXlxVHYEB     400     110v�;�RQ�Z�Vs/`-q�{�<�V��i�k�OC�C;#�SA�b��\�����r�b���ܠ:�_H��nS.�U�(G!��I~�����V���"�i��^/����S �X�� �]���2�G	�u��1&��3o���$��Y��Sz�N����.R��f����5�ׯ1o�I��k�1>D�Lʬ�^�^�����a=�@����v����l��@N��N����T��ɚ|>#]�H�[~Թ��"�x�C
g�Nk3c�`>XlxVHYEB     400     110C(>#1���Q�:������90�\%E�=����$�)8ɷ;W��B��Tu$���n_	+�HS�%D��-<O��3�*-s�N	V�^�D�U3d���Y0��0��
���Y�B!L��v�'k�h����g��jg��\O~�{<��3h�X�:�:�E����>����U�����X���B��-��I_{T���eN'l�=eua:��)��F�V����L�����d�.-����� �Љ���L��?�NX2�4;�;d�}�'�/�zɊ�XlxVHYEB     400     110��Z�͐D_�C�|�J3�K6��=���-<�F+A5�ۺa_ԲE,1a��c���It��L�`&����ѝ:s����\�Yfn�lg�Q�E����͊y:�k�s�C_X�,A�*(ο���Ưt鴬���i�+-��A�˳C_��G�E���x����~�/&�C�OO�������ɟa��,���xmi���v�W6�|�,�*���un�^���Vۻy9�i�+��3O�b'��Y�~<�nԘ��ncs95�`�[��C��,*XlxVHYEB     400     120���֍ox��j�Zi�|H�^�t��&M�Ic�$�	��1�%LI��>���+O_*�%��m��n�:���:̼�2,�����8s =��z�3���3�G���o!Ne[���F9�l�J��&o�}�=(�=]郢TK\�nQ�g���m���«֫H�4u�"̙��D��)8�[h�θ@W�@�Y�nMI8� mA投�鼕��Yބ_7�IAh+nw��! lc:�џ�i[�a�\�:��GG�G��XMw%�r7��7w����_�	c��#�#OXlxVHYEB     400      b0F�F�f�Oss�'���ly�|��*���G���� �w���!�ą���D���}J�qϤс�h�M�G������� Ϝ���\w$ln�&J�g?���hCaצ(��t{L�)uIeA������Ri�F�yb�(��^���h��_l����� i�������'?�XlxVHYEB     400     1b0�����t��#��T/]���{{n#��zHd�ɴz��l&k�ω6�+�ZZ�[�Q�g+���KՎ����1��>	��+XS )[�R��l�i���Q��Q+��-�����Df����x�ŻƂ��19�U����ʚJNZ�93��� ���H�epf�f�x�iV�ۖ;��y�y��J�f?C8����3�W����]��(3B+7���Ί`(k]Zl��,��¶�"Fc�ˑ����N�J ������?{�O�Z/��n���|>�K<����ݺ `1.��ns��c�qO��ތ.��(�����ۃ&�?��13�V� ʢn���q'�R/�⣒��]�[���\�,�#�.��rC��~�1��rjWJjS�*1V�vK��Tcy�� �Sa��K!��^2_W��ڦ�K�M�zY��%XlxVHYEB     400     1b0�C<��r�}8�s<an�����EH���%p�g�6G�%�f#^t47jE�k}�r��Z�1>��_����do/�8�r~@������8�U��L�9#����T�f��P6ZP�1�G�I���e�j���܈wp�P} ��
� �]��|t=�����G��e%(��
��(����w��Z�H�UE!j��|H��e�gQrʳ�Bób��*��`��H��z��';5��r.�e.��Lը2���f�*������؎VkB�j$�̭��~�A��<ץq�j|B&��J�X6Oϊ��5�e�㳸p����Q�y��Y��+ڤ�q�  H=��y���V��=K�
]9�y����u��� ��j�d%��m��9�ȳu��{�X�)^&D�):~�l�Ԣ����ЮV��s���Ӈ��@�j�D�91Qk�[�.U_�	XlxVHYEB     400     120�aZ�� ӷĜ4�m_^W$;�w��!�����hI�]�<7?��� #�(8�cA"�MZ�&������jv�!�nh\b�]��P]����X��Q�q���9�e����
-ޫ<o���I�4�S͌lD���M$)#���Umu�Y�i��R�#��*�!�m�Y-嚳�8�zC�|[e�7�T=#�=�Ra4b2Nhj�D$�e�e�а��ᶑ�ls���������ď�����lg���uK��+�q!�=ެ]�Au*�W?T�L��N
/��ԏL|��XlxVHYEB     400     120o�ۀ�m�����R�4�0�٧����r,W�q�N[���M��k%A��i�����"ϫ��IW6��.8�q��4w�U�"�������4V\
���:,ߒ�������a�L8�tf�a�(���i�(OE�?��%�9�^g���Y�j}���m��d���_Kp���Y�dCj���q�%�%�>��� ���J%����o�+���3��l��҃����xY-Ӏ��X8�H [0B1��R������2.���ef��&2��/W����.[��#���	9yG���XlxVHYEB     400     100�m1���g��b�88��o��d��|����"T/���j֭����f�ϑeXm����?S��ݻ�[Fc��ɏ���S�/53�¬$r����� �%�[�BE�Mi`�;P\B�`j	�LLGi�F��d�M����,��l��Z�J+Wyk��ӎa��)�� �NNҪzH�'X��˯{��]����&%MщBt��и�[�A��^hYZ>��?9��IR��'���{"����úq�h�'$XlxVHYEB     400     100��C�c�G�%B0K6X�Ω��.٧��`-�#J��Ql��P���͛Kn;���r~!F�_�b��V�Ί�5��G˅z�@�bZ w��,��-���Ű�K-�H�����s���,\'�d{�ZO���@�x�<a�b��V+z�ǲ�"�7u��ZڽJ���p�����1���}���Bj�FG����:,NZ]�<�M74�c\�~����J@�n~RTe�^�)�m��G�������/{�F�<�xY����V�XlxVHYEB     400     110�Cۏ�"c��p�r��(��Sl
��7�J֕A�ruh�o
a��c����{�&�,�sH���ڲQ9���5�nXD�	��9(�.Z�a
�Pa�u'x���n�ˮ,=`�=*O�����S�f��2���'�TƉф���T;���5MF��8>���wn��!�J`�\K@}Gx�h�n�>u��Vf�����@��v�Y�`H{���;���W�������L5�6&'2%�['���X�k�rA[�u���Ȟ�Z�J�w.ӥ���XlxVHYEB     400     130��=�����b��lc�5,NR0i�I!m�a�I�'L�5���D}��W�B6�������n"fd������]��v������`*��C��n-�A�KC)��'��"�T�������[B����ZȲ�8�!�l��>ڧ��_*�k;a���`��.��)Z6�K4��G����VL��̴}�1z�h���l��#G��	�f��m���0����c��T�ے�][����C�w]�S�,�9����.�ʑ�]�M����;3���uƵ�����U����E�t�}��jYb���QC&XlxVHYEB     400     1208���r[T>�E�C�Ɯ�	�N�4�@@:g��ŷ�x�,�!�Wt)k��bM8ߎ��Xx���$�ר��?��l���ca �ω]����O����f]|?�g��g�Y#$b+����Hgow��� �4��Eh��A�;��UCX*x�M�rڟ���ޕ)�����8��b�Y�m��UWx�ׅ�7���ME5��Mk�f�60p�Aq��	2���4�}�{��1GEn+a-+�F��b��)���:T���E����J��Մ ��C�XlxVHYEB     400     100�����lO��7"�����C����{1���JIoUЕv�P�G��2Q0���[�j�WM������3P�H�9�3�3�����F�Nb�mf��y��{�%Q����s���I�?��`��s��Ϭ3�v{�qp�6Sbl�1;�oN_Dlr�D���3���L�� �SQh6�ب)��.��|?=���"���G�538�p;��ښ��/��_Ym�F�"��~���)ξ$�L�ZP��I�ֳiȕXlxVHYEB     400     1b0�#��4|������(X�쬃S�Viv�0ʰ��Xy-������:r*�����jCƶ���J���T5��!��	��oS��ԣD_���t�g@�)r%9D� �g���@�d�U�kx�-��e*�����r�}�r<��B���NeT���C�,�8�o��e��f���c��#|{�!w�L�l��s�+/��5z��7Y�+�b��Z'����k����[���A�n��<��������UT�#v����a|���/&��+'�o>�|�ʬR�
��P$sH�K�i�x�Tt�U$���Ɋ�#�a�"Z���/�K�=�i��'xd0�ÿ&b�u��R�e-�W>?LE�e x��PpC��\,ŝ�M]����u�vΠ��3�^ds�ՇSB�u,e����j�(�b�e&㞔}�sq5����?W)��XlxVHYEB     400      f0/��+ >p����iZ��}�{?�HD�>�Q�S�~� ��v�o�n���v�Ȩ������WW�'!�L~%b�?�G�WHi�2�9l�&j���p����%�/Ǆ���=�9\���g ��:�9m,@O-�XL2Ev)��\�7�H��=�[�+X��
�s�%fM@��]e<�����}�����U���d>O�f�_�dװ��}W������$���O^88��'U��u���XlxVHYEB     400      f0M
�Ҭ^�hy@����ĵ��L�Ҫ�bee�����L+� {}�_����d5��Vz?�c�%\P���¥}[I(�l��`�0�ܣ�;��3�G�27t��*�6�.��`_|/�����T�f@p����� �7	i�a�|�E=� �Eӟ�ղ�̸I���an�[���_����@7��W?��ţ�ݜ��Ԓq�Lq|Ԣ��6j��xA�d�?��9�3�J�i�ӥ���������7'�{XlxVHYEB     400     1b0���neD��ժ��ֺ���i�ӛ0jS�+-�M��͘�
�n������y٭ZHس����cۑ-ӔEJ)��:�f|���+�-b�l}#c_��᱁S뗱d�#߈����k��+hl��X����E0��ᶘp�4�<U/��W��?b+� �|r��aUD�QeC;�R0j���w&R��
d&#*��R�^�ЦĤ�Ѣ�MF�h�o�A����J���E��X7���G(k."�,gp}?��&�#��j�J0��{.p3��z0����<��zN֭�\���۰�N���-5�� ��`�Rf���E(`�s���3�Ht�}��]��*�q=t
1O-G�"����޶֏3����O��@�_{�~�T�Y W���~�T���f����y�{
�.���,Kr>p����=e�؈�_XlxVHYEB     400     160�u|�I��t�i� ]q/�;�8f6�:�z��ٵ��#�����n8YQ�b�����6hE8T)�D-Y�D�;ToԦ����qs������l���ɞ�R$���f��/ _����Г��8�a�Is8�f�OR�<B;��=�ޖ��E���Y:�&~��)���d��^�4����7����ѳ8HIq�`vHv
��6��Su�Zk(S&�)�tz!B�͌��������D	E�#{��g����w�
G�����:�f���C&%c<vtk,��|��N�)8��*�c(�u�{�`dw���	���SA�}��p��`����b������j=E�M$q�5e��蠧����k�*�XlxVHYEB     400     140w��v��c˳��m�[}�e�預�������so@������M�Y�g�z��a����^8"b�e��\A�C���Jd���c"�G�|#]�k�`�Y���I*��9�W1����>�{��jmv�g��6s�:�,�%�-�>�CfK�En!5ū�<1:>�󂣳�Q��vT -�SwN>�����L�G��#���P+��徝h�j�і9� �����.�v\��fҌ���䶍�w�J�I�8�(*�g���dJn��$�FKɨ^�מ�-���"[�%��_��]��s����.�	�Jg]��XlxVHYEB     400     150 K�f9�){N)���񰃎��L������K�H:fs�����ւ� �;���~昔��Ϭq��{$��9yζ��'�dC����6J{�?QN�2ETn�C�xX,�ߘ�l�&�WbeݙߺI�;��6�����t��@����
�A|&��!˹`ƪ�H�����[J���ɷ^�ޱ;���[���զ�fr�ٱy� �!��W1I��|����?|-��2�*�+���������N�%у�P�<e�Fw�{�S`�O��X�Ycӷ��#F�LC�����.�)�&%�S����U�2�ʄ5�:-�N�aæ�ulN��t�:&���zqa4F���XlxVHYEB     400      e0��
�)����cS�CZ�����^FbJ���w����՛W�Z� ���,P�Ur@tǥ��6�,�hC���9�_f��X���1E���HU��4x�z��sα*��1f���JS��כ��c�}�=�R��Ĕ����B)��u��mZ����E.-G8<���EЈb�9�P�^�b��	��_�����s)����X��"s��U���|��oRf��XlxVHYEB     400      c0�+Qʮ��r�6:_2Ia�\-$u��
G�:��F��E&��f����mF���2���Vý��H�<e�mr�E}�L<h��f�6��QNVl˸�=� ��*��:�h������¤�O��;e���VS~w'v
�@"Z�m�PW)Ń���2*��_����z@���^٧�"11YH(�d��h��(���CM2XlxVHYEB     400      c0{�ژ�������<�&Ι�7cB�4_UQ��٩�s�+ A�:.;�r^z`�odꎈ��9�	�N߇6��{%����<9��s�5ŀg"���e�r����]�Pk]��j��'�����гQĦ���F���z���2��$�6�͊ P����;����;.��8C2�A�p�v'�c��;>j���f�lXlxVHYEB     400      c0��Oa�ڒ�/�q������^Y�X �5����@��Ē|D�lWs��7�jZ�W���8��d<q�m�5رdK�[=��E\bbJ��]
�^�Ԥ���&��H��T
m���
�����+��H�_3��	����u���TՄ�Y�k�zT�r������y��2����3�@矦����p�XlxVHYEB     400      c0{�ژ�������<�&Ι�7cB�4_UQ���8l�0��T	o*T�+wy9Z
��� 
׆z!��4���B慡�z��v�?Ś?���/&c�8�w��՞ g�%��͸�����"+=�;�T�K>���ᄾ�bm7�|y>m0������|�a	�WL\yUv�'�W�JɤkN	)bxh4y�����XlxVHYEB     400      c03Q��5�����pE��|��hĨ"�"n���)�t�����E�3��p�;໾�Ț�V0�\gM�J?��7Vس('���~8�E���r~��)�3"��o��{��Ζ*��Y�%ZX��t��ï-a|��KE~�U�����0O"Dpce�1�}�]n�$��j9�qG2�9��XlxVHYEB     400      c0��듵dˁ�S�CQAZr���Y�g`�+?A]Y4+j���&"��"Or��"�j�`q�8���yI�F��y�q�;R[��t�p��tD^V� p���F���姽n�WUz��� ��J[�񈮏n�O?ۂ3�eθ�а	ӎ��#�M��QR=2�ؘ,��(��%]^�	�W�Uqz�6GԌ�t�;��XlxVHYEB     400      c0p��+�}����vܰw2\�Ci��3�>Ɗ �*ujذ���q�ӓ���֨˄��U5׾g4v��g��n���� ?�k���&Nz���%.6��l͖�r�r*���c^t�[�2���C�L��C�Y'�
^��?|b�[�.���W�ODְD�Q��K�Q2DP8ȚY�[�"b~ҥ�qz��b�����w�9fXlxVHYEB     400      c0e`�r1����Y5F�����?e{�\�99�6�fO'n��UC��r/��������<�a�0��Ov�$��ޛM��v��|�\��
�$T/l�P:h	�"Ƅ�r>?�!$���� �2�b����þ��A;��b|��R���_�[#�<}Ŋ��nH=Z�x�-�VL��}�Vs*󷳭�)%3��F����XlxVHYEB     400      c0�o����!fуO������1���HMd���^^���G��R�:���D����3?|�WO����0��,Ǳn�f�^��O�:mtԓ�K3��'"��{������S�mcc�Z ���2�EU��0�)�R�߆L�W&���&f~�t.�����*p�/5:��T{�l��-=g���:��XlxVHYEB     400      c0���B�t*�?}4��((Z�8T���2�I��Fw~�dO��]��=�;��5������x���H�*�L�|�Kh� �G�N^z���m>�i��%v�wT;�E�1%4#u�
-~��P^B�f�6gV���R��m��C���Ɠ%V��Jc�6ώ
v?I�S�E=2�e}�g�a[/�o=��:��`ܱXlxVHYEB     400      c0�F�)@
;j(=���½=rR5�����!��mX����B�bؤ��s$M�hƅ��"�OB�
)�20�=I9���8�h?�M�@��I�yqA��P�$�X?yo������mE�g�J:ϸ�)]��.W�W��ԭ����c�
9�,��ni%���џ�G��L�]u#��\%LS��y�,�T��h(XlxVHYEB     400      c0̻�F��m�u_x�Taպ�!��N<� ��Q���Ȗ���b���#��N��)>�%M�e%�rɄϰC�3������do�k����lrW~���o���r�k�`� �i�T���e�ju��G�,�I�id�N��m��Y��HML�M̟�!�	�wj�z\���� ���w,���
1P�is��XlxVHYEB     400      d0~� W!����%����E��x�p�@�ҕ?��-s6�1E���t{~��tc���X�3��3��4��\W1!\�$�u��.5U�{�Ă�x����MJF�.�.R�t��B<�z��B��&����;���vq�
u��,��m�[��Ӌ��&�3n[�ü[�#El<�)��pWF��~X+@�n��9��;�>�tv
y�RcrXlxVHYEB     400     140/����k�Rs
nV�oA����w$�)�T�QY�c�Q��l-E�1u�����C,j���߅�A:�:�_���!Ud����M�j�zT�+J��JB,E���N��ac��/ppW*g��"��o�_ߑ'���Y)���Ut��VW�����:(-7���x�~ڠ8�v���z&��`��V� oz���%��Ul�<��H�~0D�8�<�&Y8�ߎk�-��	2�ձ4�e
�s�ȣpi
ޜQ��wAJ�����t�1�l�0�OĖ���nw�Z� p@�t:��85��QO�,[[I��Ѐ%Ѐ��j�禬���G�{{��=XlxVHYEB     400     160��jGlD ��w�m��������jW	-���(WJ{�E*L����Z$!�7:��JW�[!���$�0L�@����ϳ;7�%����E�s�N՟�*\�t@����D˳����D����Is��1�[�׬t"���U��M���i��L����R�����}�8ycA9u�R�^�Y���[�:�YHb�# ��9���!P3��K@3߼=
�Ayh��mV�$�J�6����ޚ�>������Ԑ��ԡ����z	��w9ޠ�A�jܫ[Ҏ���������x$u:s~Q�s#�5��>�G�F��)0���l]��dݕ+���׹ƫ�Q}�R��^�XlxVHYEB     400      e0�*@n�>�QI������4�e����aZY�K�e��z
�����q��9�^�I5Z��;�w�:�D�L�.|�z�Z�Z��\�=vh��F
ci����~<&��2�s3o���rt��}2h`%�֗Mo�OxC�줸�d���� �ڊ܏����v��,LcnmeI���ȏ�$?������B�E����,��>�꡹r�k��z�Ӟ�pXlxVHYEB     400      90:0cD�ƺ�*�aD�sIK��(���4)$ǭ����-l������?��I�����<�F3 ��|*.��_=�f{������3���f�
h5R������_K�p^��Z��؇ �q@J�Y(���0�^l$��`XlxVHYEB     400      90.B��I�w���$��YöW�]����� �Q>A�:�����VF�*�8��z<� �=�#LZ�KdE �n�ᦥ���*�99_�CH�����7*�*���Jn��t6Y�O���� g
��F�y\l�c�{b�#޷8��em�+���:XlxVHYEB     400      90�� 1��6�)H�Ů��1"i��H�<uJ�U�@��^���}횧��V��C����=(+v����3���������A���Y�#P�Fb?;�yf+�%���_��r �B�HN4��1+�B^^qP�Q3���
2RP�����1qdd�ڒ�XlxVHYEB     400     120q��Xo�g,�������Q])�8���&����gm�bq�|d�5B�'�u߈�m�;V(�)
�֣�ۤ/?K#7����}��k��杪,�
ثW�?�S`����C�T��Y@�D���zG�Vfj\fb:޲��q�s��+�ď��<�Y��ģK�ek<��?�_�A��N���!�'�6a���T���Z�,�;U �?P�s�1j&�
(�？�kN�S��!�o%�����W�k�x6�F� ���`x�$���?0�&�<�KTm;��!fd�-Zn����9^C`��p�?XlxVHYEB     3db     180� �c����'�����,�����R0�7hW=jP�%4~���X�?� ��4:�b� �	��i��ӯ�dj'�TUN�yg$�I$ܚDl�5�KM�|���M������EQI3f�j0m+��Q����<�u��VF��ʹ�@�<�~69s5�A���1?�*�y����t���CY�RV�E�WN1�W^�J�����*�JU��-� �O�:~�*�Y���{��b�	��w�������d�ᷤ^����o�;<~Q�Z��yN�R8�>�+����U'������8Bxɪwq�&3�?,���M*}
pA߲}e֋�(m >�jpQ��V�`A��l�.��ʽh:$�XĔ#2��8d�D`��/���b�y�6@�� [�