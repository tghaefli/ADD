XlxV62EB    82eb    1650�d����lt�G�����Ԍ��/�b�aj�.��\����W�+�\+R�8�"Xh��q�c'�V�G�,��=~"=D���$���OC}ިq@��1��A��r߁wQ�䆌S,��h�g,��D����v-?�	?�_M=�Ǔ����ݔ�.?�I*]8��2a�� �����r�J[��+!�f��)l�| �7�u8�ti��,���]���q/���e� �����Y����@f2A$������i������.M]�i�S���#����ӗC��;��j,r��m|�����U�� �G$��*-�8�n9��Ν�D �z�N ��gK�mV�@g��Rǝ��֫1���ͩ��n�����	bDK�9]�R�֋R`�]�9�;�u���5�����p�|w4�QcIl��������]�[)'u�UWZ����� s4AT�(�D�A� ��Dn��8yx؄`+$��H?L�ԍXN7�YR�`K��6yC� +աm*G�\=�d:�mq5�iRV��P�ӡu=��Xcڝ�*�8i��Z�2e�� �x>�xQ<`�I.
N[�	�ÞO�Ng�%���.#ʂ�w���7�
�	�o�#ﰔ��7b�et�T�Qq}E���{�=�9,�/Ť^�r�G㾎��y8l6�w�����B���^a��L?1�M�5�`ǅQ��~��U��k��i�Zu�ʇ_��$�'ַ���j�/�Pɍ���=o�@���z2��>{�SL��ҽR���u7��B�Q��";�؝	Q�HF	U$�a�BTmϡ���Ũ��M�`�&�v���v�bC��	C�N�%�M�M�/�M�a�K�{�˞��L�s��m�siG�L�����^��?v�Cx�;���Q�x3�w���v��4�W�in���v��5��W��zB�fR��Ok�@�
�W����Dؑ+��s�E.y�g�H%?����Ҥ�;�P���ܭҞ����4� B������P\=ݹtN1�.���Kҕ@>m3$6���Q�������-p����\�Ӊ�hĲ 92����H%,/z�v�t>�s9�M7��Po����˝Y���G{�� ߬��Y�K���{�o��Ld����D�Я�W�kLb��~\ OD�����A^�k���'���aB+�(���u��D"f����������
=��u}�"����)���nS��f+�������fâH�K�o�B�l��r�H&(9S��>Tކow��*����fB�!w�/�>����cp��b*���-� "x���֊����9h祈u�ꤙA�6�\w����P�;�~��KY�5����=wh�u�ow�e]�0�ɻ:eʠE�y8e�:�/�х~�G�Em��hl��$�:���;�2�q ��$����唩��f#�A#B��7�v`� !f���H�s]��*�Μ���K����n��G�	.w14$�	�����5�,�t��`����^��Õ9�W5���)0=L��Qi�����Z�_jbo+k�� -7s�Z>��ē+�5����ۉKz��&��u\���*��� ��y����?s����rٛhU�fT@������"7�����a��9���RƁ�k��c.�+2g<	/��@Mj�=��iw����I:E�%��G+k�JjY�Z���O_Yì���w1v��X��3��P��OT�.��RAW�	�'!���^,ӓ��"�Ψ����)���R�������{
�F[�)�"<�cB�Tyx�6�B�1�(`�O���.�R~Ą,��V�T~���xl��n?�ShҒM���˴�c\�yy���@Μ��^�4�oS{{B�"�� ��՞Y-�Qɼԧ@d�'y�/�[�1[�d��m��4�	�����ƃ�f[�������U�t���Ou�ǣ�,zpU�G0� 
�e`)<\H�S�z�e7J��QUE�����H�PBպ� �"�0�:�"XI�n�k'�@S!���D�SuSVQ�:5���2� ��?u�a�}f`$|���ӯ���$?$����X k3tٮ�sK�/W=>[�^"��ztg�';�����d>=H��+�>�1L!L$�S;d1�V1��{<��8�8\8����LU|�[���.���1H!�I�@@��h�O����WuوTI�K/��̈́���nM^j��.� z~"m��$��Ε��z������&�]�"U�ϐ�xj�4�:6s��g����Wjߩ&7-u.�o&I}r����II��=H�����׽t�r ��G�OC��t��#���i����00{���I���7���(C��L;+g�:�׀7��G�n�^�G)�A��=�ȵp�Է8���c4���f�_?[HQ����,z�cݛu��dz8�`2����v�Q�����©�����Z�PS�4��˄@>B�툆ÚY~�_#m!�H�?�D=�̾�Jde��AFi�!W @���&��O~�L��ф����aK��/�L �J��q��%R�5�� ��	Q�R�O�@��)A��e�(瀧y�Ze���
��]���xz�Տ5B�"%I������Rc#b7�xkp	7�c���G�~|��5�dl_ ŝ�疄�\�?+��r���l*�ﺏܤ��C�=�?�Ja���+�=�u.G��'�}���v�<��<���W?�o>��͛�[�8�o�C&������* Y���
�nsW��C;���-d��Y��A�(��QY�j���a��#��9��h��?�`���B�!�2�y�U����>v�rG{]�,�/���aE����4���Şl-lt{p[�R�;���Q �G��.���(/e�L(F�H��z�}��j�̘9n*4���Eݿ����V��.�r.N��w�Mm��K|呻V�Q�)ml����W1/f��eu�:s���{�!�&\�k����"6��@d�,�ַϪS�K3tꝡ�Z�ř&�?;4;�����t�$s�!�О�A옽�$nh��2b%�N[�?wmR�ܛ(ٲ��n_�/T�&uQ@��Vd'�cua�hZ��nFЫ�����,�WO�߄[��f��o�+2��%B4�5��ڝ�R�t®��?V}�[s�M޾���LGZc�!�GS�KH��U�\[�
H���9�`�93k�DH�X&��Zs�Z����Y4�B�.x�y������OF�e��M�Z��3�N��zچ&����H�LX�� �5�ىu��|���
&K<$p�������Ѱ׮X���l�G�~��+<��	q,!�187A}d��{���\|J��%'��Ar���%����t Hw�z{Raq��UKL> ��.a���'����(I{�X�><�P'�/�Q�e}��оZ��uׇ!s������/Q/�P�̲��H�/>;��7l�ί��H��ׯf�_���;�=-&ɐ<~q��/?��p�q9�&�c���*��Cd]t�}�js����5�j�Q��.�BV]9��fL�_��Jk�C���&@2�P����������%W���~�$+>A������5s�L?D��E�X��"�S���E�f�6���r?�hl.�D�9{2}��a�Nࢾ̶�>�����ݨ���[o�OX�׵��n�sϭ��������(��|��kS�LI���`��1��pf!���cܛ�R�`�?o)��+e9%��=��D��jYrɰh� ��+C���ˣ��H�cð}�ٿp��p6SNB�>'m�=^�׹��X�lJ�@��\l��$
����8(\��V��,�*���Tk]����;�>7� �]�۟���U�W�1s=<LH&�m�J�\��kE����S�/���?vm��idEv��qd9��a��s��m,��9����@����j�u����,�a�İ���.�4�w$!|�V'Y�zt#�{v��G��w:�*�P����_�O�%2��ꍣ�>�e�'���1�7%�VD���v2
���`?�d�<�����T�P���R�Y����h�4J��UY�GBQ[ڵ�v͠l�`o�i�Q���k�3��l�J�����j�A�a)�������O�h�)e��86�c��?tB�q:�,al%pC����pe:�2/a7qZ0��@$�b0]j����.��b�������������Œo�P0�z?n�ς�eu��:���^m��)���ȄVQ�P��|��벑��t-U3��-�l��z�[��y���z��TQ��\'ꔋ61��	�1�yP�?��2��]���|���]��(
~�����㌟� �^�I�y[�d�ϻY4E���X������T4�K��yʨFU4�g��s�<��k|�Zx/i嶫��"������~��`B,ݨZ�T�IBBCD�^�X�O<"== ri�6���� ����ޜ+*ӭ�a��&��x$�����#nδ)B��3ߎ�-h}�<�Ӝ��fg�@d���ݢ�l�L����rj�Ud��H��-�b�_�`~�F�Ry(���7� y�T8R���Q���#j�r|���ߏ�&F�8��:x�8V�잿�_f�S��%�[�l�"d8q���JF����g/�p��OW��I�o��nͷ&�sL�U�只�tި�	�hp̨�JZ��]}��,�c���R��,��D��IN�"����#�sf��mxY?,��Ʋ�n�CU��b��{�/�����=�Q+X�"u� �l���j	oZ9>�vئ_pg~� ɺV+O�C#^A���p�pg�8IH�w�1ttF���;O �`���:�v{,��a%:J������+]��@L��"Z-H���Ȫ���%YP�/Nޜ����IBŉx���u	�z�ƛ���M-#�QƇ7��)�b�m��q'9g̸pƇJbر(0�QcJ�ݟO�2��+>�����/9��6�C����d���7gԶ��V&��ל�[���{����߶6�S�>�s��h����9�v��i^���,~_Q,hK��������Q��(�u���{��y�͕KQ����C�6����S���&@K]e���5�t-3�e�t�)I7ną'p��
UR�-6]� `!D蹚�g��ф�o�fS;�C�b�C�	�����v�\�y1�πYF\���/��n9������t5��9�e��e���5+��0+��'�y9�d��{gD�P�c����P�j�93(��!�����*�� ����~���Uɔ~\!^M=�MS�MQ@88�W��
�.�BR/��jӈ뮕��u�P9x�>S�� Ԕ#q3��"�yf�z�M�+?���I�M�B�Я�G�=�ä�`�&Զ�{��X��Z�T�˖��^N�^��"7z~�
�n�l�枪�/���4��jr��{�N*�v��Y��K��ꬭ4��� Q���avo
�	AN�LT��Oh���mJ/"7$4�T(X��ߑJF�U&<%���U�E֖��k[�W�7MR�g�q�3�A{6�+��nR�i� �Cs;U@b������b+�2<){��L�1�Giq�q��:#���x(���y��՚^]�2�o�u��@�_1����%C�c�%�����:RF*�QV�*8�M�"