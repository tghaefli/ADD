XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ݩ��1Y�@a~������<�@�;u�ڀ����{B7�37|p{�=��B�hN5�WD�{N	��Y�*�m2��;u��-��7�#��G�}���[�`��33RV�rU��Np�&�n'�h��n��<-k
�;����y���3��(o�o-f�L�ml,�
Ӭ�X_Y��cw�I T=ȾR/���԰5�BKG���f�z$�J[^mm�޸��	Ba����A>Q����#����@��B�˵����Z6� .�;�e�?+r�Zt;F���em����+�-�a�~!��KA� d!���)o��l��/1�1x��TE�,x���}g�����Ma܀;(�-�ǔ���7�������?;���]9�9R1R��Ƕ��87
!�ZgSrd�3�:�՛�h���m@'��Gi:�J	�_E6�xld���������# �D;}<u��(�Av3�M�4Es������^�I�6����8�QL�����2qC5���1͛e�X����1�0S��O;�<򊬎�K�ˏ�m�KY1ů��$Hn�!G�r�Q_��8�@�yFպ��+��yK�� ,PTu0�t��hn��|L��K�Py��d��5Ĉ�n`кk�I䎙p�Ϥ�(NW��2r��u~����e��!{r�������_��H��
p�K�$��(��������nhF^�7n����&�,�=��g�A־�m&�4��D-�PV�+�`������\�a����`�1�6COXlxVHYEB     400     190��E�q�����kK�9V���Q,x;��?�&s�5�zxW��U���}��'��'̅H
�^E�#YW�w��0ֺʻ�٦��t�ȟ� ?2E5�R�	A23@F�@1�rq���EQY��g�6�L�n�2�iNv��;f��^��f�;ґ�Iw�C�ؤ�2u�Oi.G�ar����2��ѼXm|���<*}8ԼaQ��Sn��p*R>�� G�CI����"N9Rkm�8���;)�Ԗ�Tp��W�W=�s  �Hk]u;v�z}�! �>�&��1�4�"~	�w#e����P�"݁�$D��ٛA�>饮T��'�,���0)FL ��"4&��Ho|����@�oi��ȷ�7���6ՕR�>R�%�ݩ�q����GK��XlxVHYEB     400     180��O0��ii$ʴ׎"5[��eŒ�����'��P��ui�*�7�e�H��a�]S���K��Ȼ���>ճJ�op�%H�����) �t�1��>�R��{�ü�b3�U�S2w���M.�I��s����ݵ���Y��ct̢cgoύ!̛�i�h4X-�C�pYN�x�z?w&�_� S]�Jc����0��&�8gtA@h�"�^e?̌�U6��wCʿ���@1�U�˴��嶗-�	/�6ҎnSjgҰT�8��uF)����T���K�R ��I_J=}L�e`�:�rmT����X�H]p'n~�����a5#�]��2W�s{�'HH�,����Ik�<��"��,Q���)�f�m ��j�v���mZ��:(���g'���XlxVHYEB     400     190�B��!���&Lj)�?���g�����R�~cHz�����JQN	!a:Q9��i��2��-���,8��N��%=v0�� �Z� 4��G��R�����r���¶�����5���!��ܻed ���N�t����#�>a{���aB{o/A��*(��Ѫ��B����=h�w,CP����oj��.?�8}�f�M���"P|U�5 �������&��?3�k?8꽝y dڋ+���q��=�9z���W	�����pE�¨�q��S@��w�[�aA���v�Y���1Ȕ�u�q��V��=������@��>�Ǘl�i�SG�+%�}���DC�^H�[Iٙk�ˁ1l,#0�"����*�P�IB������t�آ����c�r?�XlxVHYEB     400     170��x�剑m
�<�o�z��t�D���0��Y�*]�8����aS0	1�Χk]HU��G�#]Y����^*<�8G���b�V��,j�TI�� J)���-	5���R����x �߭H�i%u�u��H�0�����~�j�}h�U��<% ��؈\����"y
r4���J�+�`[$�5�Et&�wX��>`Ս�G^|�?�F��=2����D�(��)�3?�/}o\%�w͟e��@|0r����d�RnuN�x��Up��)��t|��v�O��� �M�s*�Nz`E����]�K�#
t�ef䑇:��3�j�^mM:�j��B��v�~0�������	�:5*���p9��֨�	$ѡ`5S�Z��]2XlxVHYEB     400     180�|+�H��d'%
���H�ot�."���7�vQґ�0*2p[�	����u2иȥ��\-��	L����+*qZ�"~��y��|��#�4H�i7�!&7�ze��7]�D�f��IM!�{� �U�m�Ñ��32�`m(�a�ow���!C��q����M��ҙ�ϐe��Dh)�\�XY�.q��`զH�h�fǵ�����Q�^��9K4�J���?2���7�qr�v<�_IC��O7��6�bXm�&�憚��cj��ɐ}<��tĺ Ȁ�� ��[:&E��Q#���"������?��CM b�B�;N�8{"��=�b+���O�FX;����V��W�V�J��\��ڝ.�{e�~R��z�e�l+XlxVHYEB     400     140���:O!�4��DG���D��V�b1�M�Rϑ$~��*�;֟M�K�]iW��	�bQ�e��ԫ_�5U#M��xx�tX�|ݤ��Pඖ����t����R�K�U��~��a��챐p
�u�5?\U>谽)����~�ŗ�(٧�4��o��S@���vY!ߥ^#$F��Sc-x��:��)������!txG�b���X��v�E�k�؊�?�j�e��G���l@�t���)P��7��0k�.��j���_"��l3��\�l��-W',�Q�?�}�\���!��B�ni?8�H�NJ����2�!LA�����FJ�
�XlxVHYEB     400     120K$�ZRؙP�2L�@u{�����r��F	�\"��12E
"�o,���"�'�D�Z���d?���M�%�A9���f�)};�y�_����wNwI�^?ҹ ��Eٖ,�TaAQ}Y�1C���&u��;�ݚ�<�]�Hz�v�{�=>�U��9�.��M�4陙z����&�!&�U�?��m!h���� zd`����J�W��;�C	��D�)q(mU�%�Ϥn�!���Y�ϯB�HL�=pVԇ�K�x��-���xe�X��O*b�><a^-3���1XlxVHYEB     400     140���5��#G�1 �5f꘣)�����=LLD��mV=�ƈ#���$��fm7~��z�U����vW�ը<�>��G��aJ�Ѹ?b�u�����鈟�f��1��iApb�t43(��Jr��	��8A5m��3�d
)ၹ��W ҭ��i"6j���yF��4�Q�h��N���}V\�f�� �ο��E]U\;�h�o���bJ&�D��X=	]*�Ӂ� Шz����ŷ��9�N��J @�`c?�s�^��Қ� Qd�NF�1�72~l�ʘ,S��Ys�9�ނD���.9���WP��*c�.A��6����|"XlxVHYEB     400     180iY�̱���_�R}7Q��@��6�z��W��$�_qǬO�q�$kёA�W��׷�r(�q?U�f���g�@/�W Ț��:LvU�1�y�Y��T��3��bx򏶜?F� ��S$gO^�9���>�do���R���dV��L��;�@b1��{��e�.�Df���S�fMZ!��z*���h�x�����=Yi��/�rp��y��PxaȤ�{�Z�ڞ��	8�����o����P���,���k�"N0q{�����Q�5�X/|��՚Ծ��æ��I
�>T�L�WK��=?�BV��w���Y��J�7�7Z�����y�L��tHb�j$}��RCf0�1���g�y��gf��[�E_���e�S�IE�XlxVHYEB     400     150R:l	ܗU�O��=J�M����S�i���G�$�Ԙ�hP�;��a;G��a+�W�T��p���}��ͪ�ٺߩu� O1���� G((���W͟f���>
P�g��������B���佢�>�9���@hܫS<�bY��7b=�we8��{Ԟ�x�Uu��� ���r8i�"5d4�w������A'�H��z��>��a����L��>s[3�6G9���|�){�#�G7�I�Ԭμ:$SL���"u�q�:8�!=���CXĊώ;?�w0I����+�8�5�\y���e��I�O�yU�]F�/.�Ҽ�l�+��ҘXlxVHYEB     400      a0����+*B�x����i�ߘ���)�$C�>���N� S�ܗ��6^�?�AI��tÿ%57R��ҫ&�S$L�[|.�Q��H�I!��[+6�(O�W��?�a�`Nk3W[Ut�	�2�>��ZJIn�3�����c U�Vm�?��s�k����XZ��XlxVHYEB     400      e0b3��~8]:�d#B;�)G����ݫ,k\��J7�
)C)�[��� �T"c���Y����|ǈ���b�'Y��_��>+AĆi.%5n���C4��~����R�ɨ�!��jw�������Ws�H�FCwoh�\4���q0e@}D*
w��^��"@)�$jK
E�-�|ۈ��33���2O�ֿzh�]��U��T��V�h)��td�O��Յ,(XlxVHYEB     400     110ZZ`p�ٻ���9��4��H���^��	'5kqq	``��;G�hq�M�
v$���g
e�rA� H�L�u������=�v��K��;�5�2��._���9ӥB��Y*�o;�AY�J�6Ƶ0I�	���F�+d����۝{����@��qӔ�Y/�Zn����-4�_��R��9h0I�|.���%F��Vkq7M8)���%�v�W�i����=|��u�彩�C����zC0�d�ʹ:^<7�6�ר��0m����q9�#��;XlxVHYEB     400     120�G�����u'f\��3���菳&�=�j�ȓ��?u��n������Ss�����; �l���^�����n�"�9��1�%у#��v�eDA���A�Ċ��O�L��KM~[�T�lv|�z��`~J2�Z��B�h���&�?�ճg5�/ v��Jv���S��>gX�n�{��+����<V|���*�Z~��Q!*۩s-Ư�7�u\��$��(=�AS���?�����%Ѫ�a!M��.a�n�0R��S��: �R( ����A�b��~Ow/�HJc�TI���GXlxVHYEB     400     110�����i�0��5�78�2DN���ʂk�H#����N1+E(H4k�4H��n ��M8E�I�o���ޝ��؅����++���K�"�c	(X�÷��ܱe�*�Nю�ng?/#k��Ȍqٽ�9.rb|�۲Πr�5}�D$򃂋V��&��#C�^f�� ��y�t���t�k�J-�`��Vo�S�K�MJ9:j���vt�-+��N�i�J� Q����q\R]�s�O��9a��ou�1�I�V4%�QR�~�Ri��/홭MUXlxVHYEB     400     130�;��.�M�+�9�����mW�;.g�\C�C����������1x����f���LB%�sQi�|2x�e�D`�qW�H�y`-��5�U�4�A��3�~�gP�Ŕ �|^A#�@.3���Ŏ
�ړ[��p�N�(�Zߕ'rS����]���Ң�%�7�9ؐ����ɟ��^��0����춖{�gZSl�F��k��3i���¸����������T��]�]��`�����9U%�2��T��+�;X=������C���kqr����b ���R��c�XlxVHYEB     400      e0�69ٽfM��Zn���g��ZiSI�75��Q��>�r1����q�r�'���N��w� +����rS`	��\�8���a̀�-��D�Jk�8CՑCCfZX��EL��&�|�J�AE�B(�rc���:� �޹X@Ǣ����n`2ŗ]R���F�DU�\4\e.Ww1��Gx���Wk�t�ҿ.N@�K�0Q��'No��m�CJC�Ӝ(:XlxVHYEB     400      e0��,�綮������3���n���UI�i-O���(6|�ͳ�"�]��$~���H�Ue�L*�78��)�;�+�(Ƙ�$ 3��r7=z%T�aY�h���E��{��J��Iq�]즾�u)P6O U����٠�-Ԕ]�k�İ�A�����\.>�4J��{�H���vwU��bA�3&\�t &���O�(��ʀ7��'�G$OI���h����b�z6u��N�XlxVHYEB     400     180&c�	�?iy��#��R���TjX�����@3�yA\0ã��d��K�t{���z��f�X���W1�<��M��$_fD�@s��G�����u��pLU�L���7N���T��q���/0S�'�U��ݮ^/�(z�R3z|�<<�ZGK�R
��}�Σ]Pg�n���p�x��JG�ӫ�9g�B�}�⋱�%��F�o��z�v�����DP	Sҩ�6WR������`��s�2^���|�[y�1Rw�T���A��ŵ{�ߺFE��XHƣ��.B*�F�r�āE�б� @�@F��X����n�M+��\��HX��iX`F+�c�Ō�仵mkw�s��8�����*,��Kv�VpQ��d�r��XlxVHYEB     400      e0�&�돈���I3�迱��H���.��Cݍ��ى�2Q�Z�SV[�S��4  �e�1 M&�0O$��{���"���^m%uE6�o�0�gI͗\^��Zh��Q���0�E���~�6���Á{�����R.�T�!�C6�(���݇��(��*�Q��8�5ڏ���/x��ׁD����K�2K���Ӑ����1��?��+�f��f0-�����[X���XlxVHYEB     400     170Ugnօ��i��C4W�?D`"e���f�d���e�\�ogn>l�r7xFD�W-����(��-%V)N�T�����{�X�Z��J�'6�M�p�kch��j��彣f%���!$\  ��.��)�φ��e�O0 pycY/h����Fg��iB	4�9���6$��c��՞�oE����[^^H�}�t�5�<�>J���1I�>~S0��ck��V�%�@4K�������k!�L~lA��LAv��l����g�f�{�e兰Ef�+��5$̧!`!a���Wz��Pvf��X&,&D�3��BkW��>>#����'��ʈ�`�S�X�|6$��9O��k2��Q��͜H�XlxVHYEB     400     120�!kf�QE�}�z�1�);�H�`E
�6$�#���Y���Ob��z�Y���L`�X㾸�L�/K{���Dp|�2��V�t���*HqY
��7dG���'����b��z�&�BaC��B��~�ΰ�j,��l��v��:|4{�H�7`nY��x�G]2/XM��<����ج7��-[*�^�N���-����͊jV�i��m��W�Mn���7�a�RxOq)dc����gڛv�H��ڪ�b2�O��:ɪ�<�Ʒ���^�H����Xz�q87^�!F��XlxVHYEB     400     160�<a�=�]�޼�Ѳ��U��Z(�YrV(�cK���H@�,���]Y�Y>��x �.�1t]>�HY�{�rsg�l������?"�J�N��Fa�nH����!X�d����qs<X��z�RByQJ�R�j�ʜ�s�`���kgf�S�B��?@�(W3D$Y0��X:Ƭ��E���a�7�ͼ��.¡��MeL�����J�������I^~�߶Z0(�E���O���� 7�U���z��"����zB�zC��#�>��O�2��0�e�
�0�aRz��?\�a�&��lmzs�}O���r���~
+�y�賔�NҲ�{���G���DDwi�4K��zXlxVHYEB     400     150� [���1�M
�Q|�@���DR��TY� �7�7�/��Zȩ���{{(n��qsU�<��t.�"L��rލV�|8�p���ڝ�6�j��Ɋ��r])U�XA��ui�mGְ�[�j���J�QQ�����Yj�'�o؇+��}[7�@�>��қ�%��3�/����2&a �cZ9>J�QGAb4#`h8��rM��LUڹ��H%;��o)r�>��b��w3�\�p�0�n���N����ᦶ
�'�h'V�D4٥�R�Җ�Rx����G�] �o?�H���ȅ��_썽rJ_nJx�nx�kDu�w��v�}m�9?��(@
�Cp��4��{�D}��XlxVHYEB     400     1003���a��T�/�����,��6�'ô���T�h��6'�X 0{��+kF0�w�>�-�?�\r�ٚ�����d��e�*]�r�m+8���3L�I)-��n�ߛ1���kb�2t^�s9���	)�Ŋ;�����(kBD�_��(����sb�lӾ�,��=Cr"����]��X�}��������YE`*�R��f��*\MM��9.���.4>���WiiX�bK�t��Br�*-�FXlxVHYEB     400     130�,���|v��νD�3i�Y}y��-ߙF0y�/=��ᘁݚ>2���DBoZ#r��^U�&r�Ү�e��N���}>�ShE! � .�!�E��3fF�Ѹ�^��P���7�W��(����>q�F�� a����>���G�e�c<�W��&��"5�d��%��'�
۔m�E��ц�0�d1�F�;���б9z�O��Y��RJt0��l�h ��gC�^����jm�4Q�*�=������|u��h@�=W�Dg�(D�����	��}ۥ��C&\|a� �.
�=Hw_�XlxVHYEB     400     1209J�϶�3��ƃP�Oҹ��߶���=T �t0�t��eyu���dpn����[r3�8ڟ���6��hoH��i#��Y��b�=�d0�H"�#�[�TaUۃM�|�����@Pj�!��\�]����Z]�q�b_)�j�$��hYuybKj��������Z"���<�|�a÷m�Wg�C2f�K�ߣw�����i~�C�o���Z�uwڿ�`]�������\5�X�fu3����&���LV������4�$��P���8������) ����Tf�����O�XlxVHYEB     400     110�L"F�5����9`ͅNu�	2=t��Eif (
�m	�|�Z��m�$����j�F�A^bL&�z<V�^�S��ʡ�DI�J1�`���#��zK�k1��ƗBU,��|�hm����d#P�D`��氲�A�*ݔWah��۶�Ln"W?�~��=+��ld�+X�����7�s[~���D�'��W�-�[��麁�]�9��PLš�Һ����Q���4^�-���F*?@�y՛������iP����tu�|�>u�R�$U����e��wXlxVHYEB     400     120�Oޞ���"v.&��73�`
�vKKY�������o\e4Xo���X&����S�c�k�`���}b��-�M�=k���.Ւ
}&�jǋ8B�qb��v\������ƽ��V<�y��])�|�[?�.Nx1Tz��!n�����V��]�`p8��,3�q����m�e��:4����V��R �K�D0�r�����MM
F֤�Ўij ��[M�t�^���[Ɩ��� T��^/g�c��,��%�F�|r�i��x�cr,`��o\�5J)E�M���"s�XlxVHYEB     400     1c0�#�)�i�m�#���8.���Q�8W�!���꘢��F a�'פS�ٛvv���[�P5�I:�R4������4�O�l1����<e��O�1����MmU"����e�Ʋ;2��{�����H�f��c�����S���ps8^����P&�! �_Ǫ��l��,4�[!85���*zdh��e�&�1"����9�d뵚�^�`�PQ�9&����*�O��i�!�R9Q8̖��9��w����^}��;��tj�32�2$�S�S���c0#"F��ruV�&%��C�B�Ϸ��!�`�����4_e�
J�ir]K|<メ|,~�qƹ$��4�����f�[
��e#���%	!�\�o��F���N�n���R��|-�8�~�,K���q�p����z�y�P��pݕ�6g��/����spm�q:�`�,}k�68`�G_X)XlxVHYEB     400     120�Dbt����%�1"d�ԞJՏQ��3��,泗z�'��4��c����@v(ɝf��	}mG��b5��'�x��H��\�5)awE>B�����5E��������j�]e��\�=�l$K�Zl��_	S�D��Uw��i���gD*s��.�Iwk�G�s�k�Q�s@��{D���OI�ޣ���'� ���`��hCoo�,��o��
�"����߄Ƞա-���K�C�/`֨�ڻ�0j�$����\v�w�v$�:�BSXrm�l6bt;\���XlxVHYEB     400      e0P>�'Wʘj#��M7�5�Ș|Y � >T��E�������%]+��*fV�NA=<M�z����iS  �\X6��#��V���$��/p�H£��U��t�f˻��H����p��W����q����.��'�S:�8��G᧲��M��Ϧr�I�lε~X3#��QW�q����F���z�����ղӼ)�`M���߫�+��*-V��Y���
@����XlxVHYEB     400      e0��a�b�8���("�,xP
�+�5���/�&-]���Zc����Z���`�/�{�y�g�tE�ݏ��n�	�?�!�@+�1�Y��g��ʶ������z�"�vN�  � W	�T��t$��5�-���@����`U���ד6�����C�z2VʉU�3����{z(��~�j���R:�K饪�^�1X�`�qWѢ��^��W��XlxVHYEB     400     110	~t��{����p��hɎC>q���k��R��0d=�����&����H�'�(�\^
5�� v��J���!N06����c�'n���~ʶ���*��$�ګ`S��b�FF�� ������U{���4���"�������j�i#(W��_n�JΠ����c̴^�G������8��Dp��P�-:4�:�F���6�3%�jb �	��%{����7�ŏ*IzUAp�m�v�XM"�rĥ�LϮ��)1v\�5��;�Ћ��XlxVHYEB     400     150KIH�鲩?�I�	د�g�t����\"�F�-��Kw�뀫fw�f�9KG�
EG�\�M#S�O���+�7���:����JI�9���"��3��0���s'�v;���mP9חj]�tj=�-m+osQ�#ወ�l��`2��}���b:�h5���\��T]�����,���\��|���ϕ�LBT���
iĢ�*�۴B��{6^����e�z��5�.2X�M����z�fh�� ���Q�� tK������5�:�<�w ����S�K�����I�"F������?`�9��n�*G8�� c�.jE�OLr��������z#����XlxVHYEB     400     150��b�cs�yk�[��C7�*ײ|�]g"]?�`�x`�u�(G����>-(��XG�RDAHα�T�ag3 ølq�uG�iH��8���0�~����B�篘��k_���Zg1-��P���x��ˁ��PO'�E;6���j[f�t�5j7��7">z��Ivn�L� �pk�����x����[%�2�����d�1};���$kah�/h�6���0��#�.�;֯IO;�!��t��Y���H���y�a[�m�e_�7�U�㮃|z�,�$h�h.^�܉�V�}�4�֍��%���hn{�s��2?���˂��~�[���L�/��(LP�i�x�&��XlxVHYEB     400     130�_a�,�֜�
�HT�8U��g��ǖۢ�c?~h	�$gb�����̋5<I���O-I�5u|��?�e�����r�w�ً`7���ؐ��i�Qm��4�I�1�w%���D�0z��W[�F;�����C��9H��I�=��Np"���%��z@KXlM������?��1~bQ�(��L���EV[ZP�� �Fw;9
����˯m���T!���"a8����gF�e�����M�m8O��3YY����C8BMa�n�?%l�PV�q�C{��ܐJ������XlxVHYEB     400     110�\
�ĳ�㿗�Qڮ��^�&!v��d��qY_Rvp��l�p�[�������)lr��ߵ��e�H������X4�@�c�r�?����B5u��E�>�/��~]��3µ)� ;������	� ���>{�b$+��m��OK6W�5�ρ�L�Ȱt��n֍�lU�*s��^ʟ�(�O�q���\��W��UAIRZ���!M�o,��cuQ��}[н��T=�e��� @����`c�s>�*�����n�`? ���LQY1UM)XlxVHYEB     400     160�md\�U� ��zI,�=C �J/��R�@�'A��P��v2q��H��L�~O�6�!w�	0�."�y�]wl�_"���U�̀�Gc��Gvge!�����Vf��ټ��ə�^yZ��\����JJ��KP�N�x�]��Oa�܃��pX�ky7��zz�����V�<ᒴ�Zi�^������/��9��%-��2Pu|�k�/ә𪑣�6�=U`5�Jj3]�$�'��?_f��D_vq�~� VNr��SM"m%9X���"rR������vZ�&w=U)�[B[���]*5�^y�i�]�JQnD��/.|�(g�>��h�.`P^�1�#���; OO ;�ʁ�XlxVHYEB     400     150l{��	O5����"jC�c� ���d�Z	�.`�9�tm�q�WN�Ob��;wN�1�g;Px����w>�����j����NL�7B��.�p+4�'t���%�4��Y���:B�h?��_�|;m)�ױ{���	�ߺ�w�?�#7��{f��*��5�����/M��%3؃s$��߇�t����Qe���#O�H�3%��Es��du���v(��/�Ȃ}%\Eִ��9P���v� b%`J�ak�uWĻ6C�G��}�"�E�ߡ�E�"�y��Kz���nG�3��@��D`K��A�nul#��)V#y!9^�H�]��n3'��s�v�mXlxVHYEB     400     110$�6��#��t��4[(3'l	���6p��?֌;�`��)��0�I�q�O=^���师sAˣ>I7x�L?A�
&��O���9��~��"���3^��'W-�L��f`���mG'c�<~��fO���b��#�`5t�d�W���h@^���3���5Zyrh(�f5��*�,��9�L�_�$�kr��	�5��[�D�~
g?䋰Sv�_�t9�?���~�#����"� �V7i�vmv�zl��^J��E�����߽$Ʀ˼�XlxVHYEB     400     110�;�d�
$��>��xʏ��tJo;Z�4Gj��QҾ�@^2�G�,>*����p�U3'0���f��/�����lIG��Lm@c��CoB. �cC���H�EJ�����J�53?չ�y�7��l�}��2}u����
���Dք28����=>�G�i]����9��(���_e��#~#| jp��[w�fF��.�i���S�mcM��VY���>��fE���+O뇿��eT��$��ַ��={	*�f"\7jBfT��*���$�㾩R�XlxVHYEB     400     130�kz��[�d�@�r�É�����h�~t;��XU~�M5Z�qU�&��D ��>_M4��E���y|$�[2bakP����0V�A����`�b����Ҳ�\��	�����@$I�Y��Y{-Ⱥ��l�ma��Y#ϲ��6�k]��X���Q�!��Ptv�LU�|��0�`����ڼ9/0Ō���r�_LfD��\�KR�J�����bi�"5��T=A��yM�>B�[y؈�|Qj�ڥ+_B���]A6 ���62V�����e����.�.�ty�[�D�v��v�bO�s��Qm�!�u`XlxVHYEB     400     120r08��3�jǝ�l����_�qY�
F�S<F�X;~UQ� ���)�X�re ����l�X�©�^I���o��9���B�r��jȪ�X!�n���Y�D��(�� Z�M�`���Uu�4r���,���_r�yֻ~�ػ���`��Ň�a����>���dd�?H���������_�p:�[P�5Е��������t�����1d�f�n\�fF]�cy�w�
\�f�`�K�+T�jB|t'��;����r󅣍�Y�̱�}�����r%���L���ۆ$XlxVHYEB     190      b0*S���B�[y��H�e���䃾�1l��O�Gk��/���\۽��j�,M�.��+Ҁ�!��q��T8*?�:C��]>�5���ͣd�Gq0\�TN�
��<��X�&T��C�O�dŊZ��?�������?�Fv�FȆ��}�ڡ���6琢{lA��ؔ[��t�h0�!eqv�_4g��